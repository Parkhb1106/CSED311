module not_gate (input A,    // input
            output B);  // output

  assign B = ~A;

endmodule
