module and_gate (input A,    // input
            input B,    // input
            output C);  // output

    assign C = A & B;

endmodule
